`timescale 1ns / 1ps

module ROM (input [5:0] addr, output [33:0] data_out);

reg [33:0] mem [0:63];
assign data_out = mem[addr];

initial begin
    mem[0] = 34'b0000000000001100000111110100000000;
    mem[1] = 34'b0000000000011100000001111000000000;
    mem[2] = 34'b0000000000101100001100100100000000;
    mem[3] = 34'b0000000110101001100000000000000000;
    mem[4] = 34'b0000001010111001110000000000000000;
    mem[5] = 34'b1010101111001000000000000000000000;
    mem[6] = 34'b1100000000111010000000000010111011;
end

endmodule
